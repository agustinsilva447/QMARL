version https://git-lfs.github.com/spec/v1
oid sha256:d8ef30923ec5215137139870c277f740cb899104bd4b123bd391335c512235e3
size 7614
