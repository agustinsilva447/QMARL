version https://git-lfs.github.com/spec/v1
oid sha256:7765f9028c95ca5a503f7deb6c1908009dc3a47e9591dade73865f356a322443
size 1200
