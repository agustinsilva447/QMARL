version https://git-lfs.github.com/spec/v1
oid sha256:2a2ebffed5a90014ee65e3ac32fc9d9c749511bfdc7440837a2c46ad54c4d5e8
size 772
