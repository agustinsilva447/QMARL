version https://git-lfs.github.com/spec/v1
oid sha256:29d6b84aa52a1142151d7425d85466033b617b57d1ddb854f7d4641e2a208770
size 7935
