version https://git-lfs.github.com/spec/v1
oid sha256:21e69cc701acc968e8cd0018162d11277a0c867b3d973c95b1717fffdc31e311
size 1751
