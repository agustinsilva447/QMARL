version https://git-lfs.github.com/spec/v1
oid sha256:ff546f3f5c3b530de8e33b325b7c76ec03be22d4ce318092a1f72651af75f243
size 2821
