version https://git-lfs.github.com/spec/v1
oid sha256:ff9d989272181e521b7aebbbdef8e75b208a695e79225a43114482bc0be85ab7
size 4742
