version https://git-lfs.github.com/spec/v1
oid sha256:2865ddf6badc024f7cb07779f3f829b576e21c9fd1054706a827c26c5cfabb36
size 4404
