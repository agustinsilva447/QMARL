version https://git-lfs.github.com/spec/v1
oid sha256:2b6f0af96ca1ff45198dacb59761c7fdf1a7aeb90082a7d2bfbb88102da1bdc8
size 4596
