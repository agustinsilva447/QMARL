version https://git-lfs.github.com/spec/v1
oid sha256:b0fd4239428405c71618ed188f7cb3ab947f529708ac437693fd4d31bf63c297
size 925
