version https://git-lfs.github.com/spec/v1
oid sha256:000622442c68d4f7967df459aa342d9e8a64f181ec41a3cfd3a423d66edfb4ac
size 4990
